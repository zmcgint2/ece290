CONFIGURATION myxor_struct_config OF myxor IS
   FOR struct
   END FOR;
END myxor_struct_config;