-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION xor_encode_struct_config OF xor_encode IS
   FOR struct
   END FOR;
END xor_encode_struct_config;
