-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION myxor_struct_config OF myxor IS
   FOR struct
   END FOR;
END myxor_struct_config;
