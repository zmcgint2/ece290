-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION alphabetsoup_struct_config OF alphabetsoup IS
   FOR struct
   END FOR;
END alphabetsoup_struct_config;
