-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION j1bitcomparator_struct_config OF j1bitcomparator IS
   FOR struct
   END FOR;
END j1bitcomparator_struct_config;
