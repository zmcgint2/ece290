-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION bitwise_mirror_struct_config OF bitwise_mirror IS
   FOR struct
   END FOR;
END bitwise_mirror_struct_config;
