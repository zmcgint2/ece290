-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION public_key_generator_struct_config OF public_key_generator IS
   FOR struct
   END FOR;
END public_key_generator_struct_config;
