-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION XOR_8_bit_struct_config OF XOR_8_bit IS
   FOR struct
   END FOR;
END XOR_8_bit_struct_config;
