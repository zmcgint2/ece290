-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION j21mux_struct_config OF j21mux IS
   FOR struct
   END FOR;
END j21mux_struct_config;
