-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION sr_latch_struct_config OF sr_latch IS
   FOR struct
   END FOR;
END sr_latch_struct_config;
