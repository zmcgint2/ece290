CONFIGURATION signed_2s_complement_8_bit_comparator_struct_config OF signed_2s_complement_8_bit_comparator IS
   FOR struct
   END FOR;
END signed_2s_complement_8_bit_comparator_struct_config;