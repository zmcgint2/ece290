-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION pet_srff_struct_config OF pet_srff IS
   FOR struct
   END FOR;
END pet_srff_struct_config;
