-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION dflipflop_struct_config OF dflipflop IS
   FOR struct
   END FOR;
END dflipflop_struct_config;
