-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION twotobin_struct_config OF twotobin IS
   FOR struct
   END FOR;
END twotobin_struct_config;
