-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION jceasarshift_struct_config OF jceasarshift IS
   FOR struct
   END FOR;
END jceasarshift_struct_config;
