-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION FA_struct_config OF FA IS
   FOR struct
   END FOR;
END FA_struct_config;
