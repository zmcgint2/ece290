-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION full_adder_struct_config OF full_adder IS
   FOR struct
   END FOR;
END full_adder_struct_config;
