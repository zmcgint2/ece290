-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION key_repeater_4_to_8_bit_struct_config OF key_repeater_4_to_8_bit IS
   FOR struct
   END FOR;
END key_repeater_4_to_8_bit_struct_config;
