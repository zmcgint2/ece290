-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION bustesting_struct_config OF bustesting IS
   FOR struct
   END FOR;
END bustesting_struct_config;
