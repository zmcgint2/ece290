-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION ONEFUCKINGANDGATE_struct_config OF ONEFUCKINGANDGATE IS
   FOR struct
   END FOR;
END ONEFUCKINGANDGATE_struct_config;
