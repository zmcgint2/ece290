-- Generation properties:
--   Format              : hierarchical
--   Generic mappings    : exclude
--   Leaf-level entities : direct binding
--   Regular libraries   : use library name
--   View name           : include
--   
CONFIGURATION bintotwo_struct_config OF bintotwo IS
   FOR struct
   END FOR;
END bintotwo_struct_config;
